library verilog;
use verilog.vl_types.all;
entity clkgenremastered_vlg_vec_tst is
end clkgenremastered_vlg_vec_tst;
